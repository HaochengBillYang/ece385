module reg_16 (input logic Clk, Reset, Load,
					input logic [15:0] D_in,
					output logic [15:0]D_out);

					always_ff @ (posedge Clk)
					begin
					if(Reset)
					D_out <= 16'b0;
					else if(Load)
					D_out <= D_in;
					end
endmodule
					
					