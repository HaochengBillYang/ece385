//module ADDR (input logic ADDR1MUX, SR2MUX,
 //            input logic ADDR2MUX,
	//			 input logic [15:0] PC,IR,SR2MUX_0, ALU_A,
		//		 output logic [15:0] ALU_B, MARMUX);
module placeholder ( input logic Clk,
                     output logic [15:0] MARMUX);
							assign MARMUX = 16'b0000000000000000;
							endmodule 