module wallbus(input [3:0] r0,
					input [3:0] r1,
					input [3:0] r2,
					input [3:0] r3,
					input [3:0] r4,
					input [3:0] r5,
					input [3:0] r6,
					input [3:0] r7,
					input [3:0] r8,
					input [3:0] r9,
					input [3:0] r10,
					input [3:0] r11,
					input [3:0] r12,
					input [3:0] r13,
					input [3:0] r14,
					input [3:0] r15,
					input [3:0] r16,
					input [3:0] r17,
					input [3:0] r18,
					input [3:0] r19,
					input [3:0] r20,
					input [3:0] r21,
					input [3:0] r22,
					input [3:0] r23,
					input [3:0] r24,
					input [3:0] r25,
					input [3:0] r26,
					input [3:0] r27,
					input [3:0] r28,
					input [3:0] r29,
					input [3:0] r30,
					input [3:0] r31,
					input [3:0] r32,
					input [3:0] r33,
					input [3:0] r34,
					input [3:0] r35,
					input [3:0] r36,
					input [3:0] r37,
					input [3:0] r38,
					input [3:0] r39,
					input [3:0] r40,
					input [3:0] r41,
					input [3:0] r42,
					output [3:0] r
);

assign r[3:0] = r0[3:0] | r1[3:0] | r2[3:0] | r3[3:0] | r4[3:0]| r5[3:0]| r6[3:0] | r7[3:0]| r8[3:0]| r9[3:0]
     | r10[3:0]| r11[3:0]| r12[3:0]| r13[3:0]| r14[3:0]| r15[3:0]| r16[3:0]| r17[3:0]| r18[3:0]| r19[3:0]
	  | r20[3:0]| r21[3:0]| r22[3:0]| r23[3:0]| r24[3:0]| r25[3:0]| r26[3:0]| r27[3:0]| r28[3:0]| r29[3:0]
	  | r30[3:0]| r31[3:0]| r32[3:0]| r33[3:0]| r34[3:0]| r35[3:0]| r36[3:0]| r37[3:0]| r38[3:0]| r39[3:0]
	  | r40[3:0]| r41[3:0]| r42[3:0];

endmodule

/*
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@,,,,,,,,,,,,,,,,,,,,,,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@,,,,,,,,,,,,,,,,,,,,,,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@,,,,,,,,,,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@,,,,,,,,,,,,,,,,,,,,,,,,,,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@,,,@@@,,,,,,,,,,,@@@@@@@@@@@@@@@@@@@@,,,,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@,,,,@@,,,,@@@@@@@@@@@@@@@@@@@@@@@@@@@@(,,,,,,,,,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@,,,,@@,,,,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@,,,@@@,,,,,,,@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@,,,,,@,,,,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@,,,@@,,,,,,,,,@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@,,,,,,,,,,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@,,,,,,,,@@@,,,,@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@,,,,,,,,,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@*,,&@@@@@,,,,@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@#,,@@,,,,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@,,,,@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@*,,@@,,,,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@,,,,@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@#,,@@,,,,,,,,,,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@,,,,,,,,@@@,,,,@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@,,@@@@,,,,,,,,,,,@@@@@@@@@@@@@@@@@@@@@@@@@@,,,@@,,,,@&,,,@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@,,,,,@@@@@@@@@@@@@@@@@@@@@@@,,,@@@,,,,,,,@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@,,,,,,,,,,,,,,,,,,,,,,,,,,,,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
*/
